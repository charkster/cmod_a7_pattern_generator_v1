//`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 01/06/2019 11:00:44 AM
// Design Name: 
// Module Name: pattern_gen
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////


module pattern_gen(
    input  logic        clk,
    input  logic        rst_n,
    input  logic        enable_pat_gen,
    input  logic [23:0] end_address_pat_gen,
    input  logic  [1:0] num_gpio_sel_pat_gen, // 2'b00 is 1, 2'b01 is 2, 2'b10 is 4 and 2'b11 is 8
    input  logic  [4:0] timestep_sel_pat_gen,
    input  logic        repeat_enable_pat_gen,
    output logic        pattern_active,
    output logic        pattern_done,
    output logic  [7:0] gpio_pat_gen_out,
    input  logic  [7:0] sram_data,
    output logic [18:0] sram_addr_pat_gen
    );
    
    logic        reached_final_address;
    logic        reached_final_bit_count;
    logic        enable_pat_gen_delay;
    logic        enable_pat_gen_rise_edge;
    logic [18:0] current_address;
    logic  [2:0] bit_count;
    logic [25:0] timestep_counter;
    logic [25:0] final_timestep_count;
    logic        reached_final_timestep_count;
    logic        timestep_change;
    logic        timestep_change_delay;
    logic  [7:0] gpio_mask;
    logic  [7:0] gpio_pat_gen_comb;
    logic        enable_bit_counter;
    logic        pattern_active_hold;
    
    assign reached_final_address = (current_address == end_address_pat_gen[18:0]);
    
    assign reached_final_bit_count  = ((num_gpio_sel_pat_gen ==  2'b00) && (bit_count == 3'd7)) ||
                                      ((num_gpio_sel_pat_gen ==  2'b01) && (bit_count == 3'd6)) ||
                                      ((num_gpio_sel_pat_gen ==  2'b10) && (bit_count == 3'd4)) ||
                                      ((num_gpio_sel_pat_gen ==  2'b11) && (bit_count == 3'd0));
                                      
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n) enable_pat_gen_delay <= 1'b0;
      else        enable_pat_gen_delay <= enable_pat_gen;
      
    assign enable_pat_gen_rise_edge = (enable_pat_gen && (!enable_pat_gen_delay));
    
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                                                                                      pattern_active <= 1'b0;
      else if (!enable_pat_gen && (!repeat_enable_pat_gen))                                                            pattern_active <= 1'b0;
      else if (repeat_enable_pat_gen || enable_pat_gen_rise_edge)                                                      pattern_active <= 1'b1;
      else if (reached_final_address && reached_final_bit_count && reached_final_timestep_count && enable_bit_counter) pattern_active <= 1'b0;

   always_ff @(posedge clk, negedge rst_n)
     if (~rst_n) pattern_active_hold <= 1'b0;
     else        pattern_active_hold <= pattern_active;

   always_ff @(posedge clk, negedge rst_n)
     if (~rst_n)                                           pattern_done <= 1'b0;
     else if (!enable_pat_gen && (!repeat_enable_pat_gen)) pattern_done <= 1'b0;
     else if (!pattern_active && pattern_active_hold)      pattern_done <= 1'b1;
   

    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                                                                                          current_address <= '0;
      else if ((!enable_pat_gen && (!repeat_enable_pat_gen)) || (!enable_bit_counter))                                     current_address <= '0;
      else if (!reached_final_address && reached_final_bit_count && reached_final_timestep_count)                          current_address <= current_address + 1;
      else if ( reached_final_address && reached_final_bit_count && reached_final_timestep_count && repeat_enable_pat_gen) current_address <= '0;
      
    assign sram_addr_pat_gen = current_address;

    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                                                  enable_bit_counter <= 1'b0;
      else if ((!enable_pat_gen && (!repeat_enable_pat_gen)) || (!pattern_active)) enable_bit_counter <= 1'b0;
      else if (pattern_active && reached_final_timestep_count)                     enable_bit_counter <= 1'b1;
      
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                                                                                               bit_count <= '0;
      else if ((!enable_pat_gen && (!repeat_enable_pat_gen)) || (!enable_bit_counter))                                          bit_count <= '0;
      else if (!reached_final_bit_count && reached_final_timestep_count && (num_gpio_sel_pat_gen == 2'b00))                     bit_count <= bit_count + 1;
      else if (!reached_final_bit_count && reached_final_timestep_count && (num_gpio_sel_pat_gen == 2'b01))                     bit_count <= bit_count + 2;
      else if (!reached_final_bit_count && reached_final_timestep_count && (num_gpio_sel_pat_gen == 2'b10))                     bit_count <= bit_count + 4;
      else if ( reached_final_bit_count && reached_final_timestep_count && ((!reached_final_address) || repeat_enable_pat_gen)) bit_count <= '0;
      
    always_comb
      case(timestep_sel_pat_gen)
        5'd0:    final_timestep_count = 'd1;
        5'd1:    final_timestep_count = 'd3;
        5'd2:    final_timestep_count = 'd7;
        5'd3:    final_timestep_count = 'd15;
        5'd4:    final_timestep_count = 'd31;
        5'd5:    final_timestep_count = 'd63;
        5'd6:    final_timestep_count = 'd127;
        5'd7:    final_timestep_count = 'd255;
        5'd8:    final_timestep_count = 'd511;
        5'd9:    final_timestep_count = 'd1023;
        5'd10:   final_timestep_count = 'd2047;
        5'd11:   final_timestep_count = 'd4095;
        5'd12:   final_timestep_count = 'd8191;
        5'd13:   final_timestep_count = 'd16383;
        5'd14:   final_timestep_count = 'd32767;
        5'd15:   final_timestep_count = 'd65535;
        5'd16:   final_timestep_count = 'd131071;
        5'd17:   final_timestep_count = 'd262143;
        5'd18:   final_timestep_count = 'd524287;
        5'd19:   final_timestep_count = 'd1048575;
        5'd20:   final_timestep_count = 'd2097151;
        5'd21:   final_timestep_count = 'd4194303;
        5'd22:   final_timestep_count = 'd8388607;
        5'd23:   final_timestep_count = 'd16777215;
        default: final_timestep_count = 'd16777215;
      endcase
      
    assign reached_final_timestep_count = (timestep_counter == final_timestep_count);
    
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                                                  timestep_counter <= '0;
      else if ((!enable_pat_gen && (!repeat_enable_pat_gen)) || (!pattern_active)) timestep_counter <= '0;
      else if (!reached_final_timestep_count)                                      timestep_counter <= timestep_counter + 1;
      else if ( reached_final_timestep_count)                                      timestep_counter <= '0;
      
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                            timestep_change <= 1'b0;
      else if (reached_final_timestep_count) timestep_change <= 1'b1;
      else                                   timestep_change <= 1'b0;
    
    // need to update the gpio pins after address and bit_count changes
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n) timestep_change_delay <= 1'b0;
      else        timestep_change_delay <= timestep_change && pattern_active;
      
    always_comb
      case(num_gpio_sel_pat_gen)
        2'b00: gpio_mask = 8'b0000_0001;
        2'b01: gpio_mask = 8'b0000_0011;
        2'b10: gpio_mask = 8'b0000_1111;
        2'b11: gpio_mask = 8'b1111_1111;
      endcase
      
    // LSB to MSB
//    assign gpio_pat_gen_comb = {sram_data[bit_count+7],sram_data[bit_count+6],sram_data[bit_count+5],sram_data[bit_count+4],
//                                sram_data[bit_count+3],sram_data[bit_count+2],sram_data[bit_count+1],sram_data[bit_count]};

    // MSB to LSB
    assign gpio_pat_gen_comb = {sram_data[bit_count],sram_data[1-bit_count],sram_data[2-bit_count],sram_data[3-bit_count],
                                sram_data[4-bit_count],sram_data[5-bit_count],sram_data[6-bit_count],sram_data[7-bit_count]};
      
    always_ff @(posedge clk, negedge rst_n)
      if (~rst_n)                                           gpio_pat_gen_out <= 8'b0000_0000;
      else if (!enable_pat_gen && (!repeat_enable_pat_gen)) gpio_pat_gen_out <= 8'b0000_0000;
      else if (timestep_change_delay)                       gpio_pat_gen_out <= gpio_pat_gen_comb & gpio_mask;

endmodule
